///////////////////////////////////////////////////////////////////////////////
//   ____  ____ 
//  /   /\/   /
// /___/  \  /    Vendor: Xilinx
// \   \   \/     Version : 2.7
//  \   \         Application : 7 Series FPGAs Transceivers Wizard
//  /   /         Filename : mtf7_combo_link.v
// /___/   /\     
// \   \  /  \ 
//  \___\/\___\
//
//
// Module mtf7_combo_link (a GT Wrapper)
// Generated by Xilinx 7 Series FPGAs Transceivers Wizard
// 
// 
// (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES. 


`default_nettype wire

`timescale 1ns / 1ps
`define DLY #1

//***************************** Entity Declaration ****************************

(* CORE_GENERATION_INFO = "mtf7_combo_link,gtwizard_v2_7,{protocol_file=Start_from_scratch}" *) module mtf7_combo_link #
(
    // Simulation attributes
    parameter   EXAMPLE_SIMULATION       =   0,             // Set to 1 for Simulation

    parameter   WRAPPER_SIM_GTRESET_SPEEDUP    = "FALSE"    // Set to "true" to speed up sim reset
)
(
    //_________________________________________________________________________
    //_________________________________________________________________________
    //GT0  (X0Y0)
    //____________________________CHANNEL PORTS________________________________
    //------------------------------- CPLL Ports -------------------------------
    output          GT0_CPLLFBCLKLOST_OUT,
    output          GT0_CPLLLOCK_OUT,
    input           GT0_CPLLLOCKDETCLK_IN,
    output          GT0_CPLLREFCLKLOST_OUT,
    input           GT0_CPLLRESET_IN,
    //------------------------ Channel - Clocking Ports ------------------------
    input           GT0_GTGREFCLK_IN,
    input           GT0_GTNORTHREFCLK0_IN,
    input           GT0_GTNORTHREFCLK1_IN,
    input           GT0_GTREFCLK0_IN,
    input           GT0_GTREFCLK1_IN,
    input           GT0_GTSOUTHREFCLK0_IN,
    input           GT0_GTSOUTHREFCLK1_IN,
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   GT0_DRPADDR_IN,
    input           GT0_DRPCLK_IN,
    input   [15:0]  GT0_DRPDI_IN,
    output  [15:0]  GT0_DRPDO_OUT,
    input           GT0_DRPEN_IN,
    output          GT0_DRPRDY_OUT,
    input           GT0_DRPWE_IN,
    //------------------- RX Initialization and Reset Ports --------------------
    input           GT0_RXUSERRDY_IN,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          GT0_EYESCANDATAERROR_OUT,
    //----------------------- Receive Ports - CDR Ports ------------------------
    output          GT0_RXCDRLOCK_OUT,
    //------------- Receive Ports - Comma Detection and Alignment --------------
    input           GT0_RXSLIDE_IN,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           GT0_RXUSRCLK_IN,
    input           GT0_RXUSRCLK2_IN,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [15:0]  GT0_RXDATA_OUT,
    //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
    output  [1:0]   GT0_RXDISPERR_OUT,
    output  [1:0]   GT0_RXNOTINTABLE_OUT,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           GT0_GTHRXN_IN,
    //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
    output          GT0_RXBYTEISALIGNED_OUT,
    output          GT0_RXBYTEREALIGN_OUT,
    output          GT0_RXCOMMADET_OUT,
    //------------------ Receive Ports - RX Equailizer Ports -------------------
    input           GT0_RXLPMHFHOLD_IN,
    input           GT0_RXLPMLFHOLD_IN,
    //------------- Receive Ports - RX Fabric Output Control Ports -------------
    output          GT0_RXOUTCLK_OUT,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           GT0_GTRXRESET_IN,
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    input           GT0_RXPOLARITY_IN,
    //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    output  [1:0]   GT0_RXCHARISCOMMA_OUT,
    output  [1:0]   GT0_RXCHARISK_OUT,
    //---------------------- Receive Ports -RX AFE Ports -----------------------
    input           GT0_GTHRXP_IN,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          GT0_RXRESETDONE_OUT,
    //------------------- TX Initialization and Reset Ports --------------------
    input           GT0_GTTXRESET_IN,
    input           GT0_TXUSERRDY_IN,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           GT0_TXUSRCLK_IN,
    input           GT0_TXUSRCLK2_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [31:0]  GT0_TXDATA_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GT0_GTHTXN_OUT,
    output          GT0_GTHTXP_OUT,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          GT0_TXOUTCLK_OUT,
    output          GT0_TXOUTCLKFABRIC_OUT,
    output          GT0_TXOUTCLKPCS_OUT,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          GT0_TXRESETDONE_OUT,
    //--------------- Transmit Ports - TX Polarity Control Ports ---------------
    input           GT0_TXPOLARITY_IN,
    //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    input   [3:0]   GT0_TXCHARISK_IN,


    //____________________________COMMON PORTS________________________________
    //-------------------- Common Block  - Ref Clock Ports ---------------------
    input           GT0_GTGREFCLK_COMMON_IN,
    input           GT0_GTNORTHREFCLK0_COMMON_IN,
    input           GT0_GTNORTHREFCLK1_COMMON_IN,
    input           GT0_GTREFCLK0_COMMON_IN,
    input           GT0_GTREFCLK1_COMMON_IN,
    input           GT0_GTSOUTHREFCLK0_COMMON_IN,
    input           GT0_GTSOUTHREFCLK1_COMMON_IN,
    //----------------------- Common Block - QPLL Ports ------------------------
    output          GT0_QPLLLOCK_OUT,
    input           GT0_QPLLLOCKDETCLK_IN,
    output          GT0_QPLLREFCLKLOST_OUT,
    input           GT0_QPLLRESET_IN,
    
	input [2:0] prbs_sel,
    output prbs_err,
    input rxbufreset


);
//***************************** Parameter Declarations ************************
    localparam QPLL_FBDIV_TOP =  80;

    localparam QPLL_FBDIV_IN  =  (QPLL_FBDIV_TOP == 16)  ? 10'b0000100000 : 
				(QPLL_FBDIV_TOP == 20)  ? 10'b0000110000 :
				(QPLL_FBDIV_TOP == 32)  ? 10'b0001100000 :
				(QPLL_FBDIV_TOP == 40)  ? 10'b0010000000 :
				(QPLL_FBDIV_TOP == 64)  ? 10'b0011100000 :
				(QPLL_FBDIV_TOP == 66)  ? 10'b0101000000 :
				(QPLL_FBDIV_TOP == 80)  ? 10'b0100100000 :
				(QPLL_FBDIV_TOP == 100) ? 10'b0101110000 : 10'b0000000000;

   localparam QPLL_FBDIV_RATIO = (QPLL_FBDIV_TOP == 16)  ? 1'b1 : 
				(QPLL_FBDIV_TOP == 20)  ? 1'b1 :
				(QPLL_FBDIV_TOP == 32)  ? 1'b1 :
				(QPLL_FBDIV_TOP == 40)  ? 1'b1 :
				(QPLL_FBDIV_TOP == 64)  ? 1'b1 :
				(QPLL_FBDIV_TOP == 66)  ? 1'b0 :
				(QPLL_FBDIV_TOP == 80)  ? 1'b1 :
				(QPLL_FBDIV_TOP == 100) ? 1'b1 : 1'b1;

//***************************** Wire Declarations *****************************

    // ground and vcc signals
    wire            tied_to_ground_i;
    wire    [63:0]  tied_to_ground_vec_i;
    wire            tied_to_vcc_i;
    wire    [63:0]  tied_to_vcc_vec_i;
    
    wire            gt0_qplloutclk_i;
    wire            gt0_qplloutrefclk_i;

    wire            gt0_qpllclk_i;
    wire            gt0_qpllrefclk_i;
         
//********************************* Main Body of Code**************************

    assign tied_to_ground_i             = 1'b0;
    assign tied_to_ground_vec_i         = 64'h0000000000000000;
    assign tied_to_vcc_i                = 1'b1;
    assign tied_to_vcc_vec_i            = 64'hffffffffffffffff;


    assign  gt0_qpllclk_i    = gt0_qplloutclk_i;  
    assign  gt0_qpllrefclk_i = gt0_qplloutrefclk_i; 
      
     
 

//------------------------- GT Instances  -------------------------------
    //_________________________________________________________________________
    //_________________________________________________________________________
    //GT0  (X0Y0)
    mtf7_combo_link_GT #
    (
        // Simulation attributes
        .GT_SIM_GTRESET_SPEEDUP   ("FALSE"),
        .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
        .TXSYNC_OVRD_IN           (1'b0),
        .TXSYNC_MULTILANE_IN      (1'b0) 
    )
    gt0_mtf7_combo_link_i
    (
        //------------------------------- CPLL Ports -------------------------------
        .CPLLFBCLKLOST_OUT              (GT0_CPLLFBCLKLOST_OUT),
        .CPLLLOCK_OUT                   (GT0_CPLLLOCK_OUT),
        .CPLLLOCKDETCLK_IN              (GT0_CPLLLOCKDETCLK_IN),
        .CPLLREFCLKLOST_OUT             (GT0_CPLLREFCLKLOST_OUT),
        .CPLLRESET_IN                   (GT0_CPLLRESET_IN),
        //------------------------ Channel - Clocking Ports ------------------------
        .GTGREFCLK_IN                   (GT0_GTGREFCLK_IN),
        .GTNORTHREFCLK0_IN              (GT0_GTNORTHREFCLK0_IN),
        .GTNORTHREFCLK1_IN              (GT0_GTNORTHREFCLK1_IN),
        .GTREFCLK0_IN                   (GT0_GTREFCLK0_IN),
        .GTREFCLK1_IN                   (GT0_GTREFCLK1_IN),
        .GTSOUTHREFCLK0_IN              (GT0_GTSOUTHREFCLK0_IN),
        .GTSOUTHREFCLK1_IN              (GT0_GTSOUTHREFCLK1_IN),
        //-------------------------- Channel - DRP Ports  --------------------------
        .DRPADDR_IN                     (GT0_DRPADDR_IN),
        .DRPCLK_IN                      (GT0_DRPCLK_IN),
        .DRPDI_IN                       (GT0_DRPDI_IN),
        .DRPDO_OUT                      (GT0_DRPDO_OUT),
        .DRPEN_IN                       (GT0_DRPEN_IN),
        .DRPRDY_OUT                     (GT0_DRPRDY_OUT),
        .DRPWE_IN                       (GT0_DRPWE_IN),
        //----------------------------- Clocking Ports -----------------------------
        .QPLLCLK_IN                     (gt0_qpllclk_i),
        .QPLLREFCLK_IN                  (gt0_qpllrefclk_i),
        //------------------- RX Initialization and Reset Ports --------------------
        .RXUSERRDY_IN                   (GT0_RXUSERRDY_IN),
        //------------------------ RX Margin Analysis Ports ------------------------
        .EYESCANDATAERROR_OUT           (GT0_EYESCANDATAERROR_OUT),
        //----------------------- Receive Ports - CDR Ports ------------------------
        .RXCDRLOCK_OUT                  (GT0_RXCDRLOCK_OUT),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .RXSLIDE_IN                     (GT0_RXSLIDE_IN),
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .RXUSRCLK_IN                    (GT0_RXUSRCLK_IN),
        .RXUSRCLK2_IN                   (GT0_RXUSRCLK2_IN),
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .RXDATA_OUT                     (GT0_RXDATA_OUT),
        //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
        .RXDISPERR_OUT                  (GT0_RXDISPERR_OUT),
        .RXNOTINTABLE_OUT               (GT0_RXNOTINTABLE_OUT),
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .GTHRXN_IN                      (GT0_GTHRXN_IN),
        //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
        .RXBYTEISALIGNED_OUT            (GT0_RXBYTEISALIGNED_OUT),
        .RXBYTEREALIGN_OUT              (GT0_RXBYTEREALIGN_OUT),
        .RXCOMMADET_OUT                 (GT0_RXCOMMADET_OUT),
        //------------------ Receive Ports - RX Equailizer Ports -------------------
        .RXLPMHFHOLD_IN                 (GT0_RXLPMHFHOLD_IN),
        .RXLPMLFHOLD_IN                 (GT0_RXLPMLFHOLD_IN),
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .RXOUTCLK_OUT                   (GT0_RXOUTCLK_OUT),
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .GTRXRESET_IN                   (GT0_GTRXRESET_IN),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .RXPOLARITY_IN                  (GT0_RXPOLARITY_IN),
        //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        .RXCHARISCOMMA_OUT              (GT0_RXCHARISCOMMA_OUT),
        .RXCHARISK_OUT                  (GT0_RXCHARISK_OUT),
        //---------------------- Receive Ports -RX AFE Ports -----------------------
        .GTHRXP_IN                      (GT0_GTHRXP_IN),
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .RXRESETDONE_OUT                (GT0_RXRESETDONE_OUT),
        //------------------- TX Initialization and Reset Ports --------------------
        .GTTXRESET_IN                   (GT0_GTTXRESET_IN),
        .TXUSERRDY_IN                   (GT0_TXUSERRDY_IN),
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .TXUSRCLK_IN                    (GT0_TXUSRCLK_IN),
        .TXUSRCLK2_IN                   (GT0_TXUSRCLK2_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .TXDATA_IN                      (GT0_TXDATA_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GTHTXN_OUT                     (GT0_GTHTXN_OUT),
        .GTHTXP_OUT                     (GT0_GTHTXP_OUT),
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .TXOUTCLK_OUT                   (GT0_TXOUTCLK_OUT),
        .TXOUTCLKFABRIC_OUT             (GT0_TXOUTCLKFABRIC_OUT),
        .TXOUTCLKPCS_OUT                (GT0_TXOUTCLKPCS_OUT),
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .TXRESETDONE_OUT                (GT0_TXRESETDONE_OUT),
        //--------------- Transmit Ports - TX Polarity Control Ports ---------------
        .TXPOLARITY_IN                  (GT0_TXPOLARITY_IN),
        //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        .TXCHARISK_IN                   (GT0_TXCHARISK_IN),
        
        .prbs_sel (prbs_sel),
        .prbs_err (prbs_err),
        .rxbufreset (rxbufreset)
        

    );


    //_________________________________________________________________________
    //_________________________________________________________________________
    //_________________________GTHE2_COMMON____________________________________

    GTHE2_COMMON #
    (
            // Simulation attributes
            .SIM_RESET_SPEEDUP   ("FALSE"),
            .SIM_QPLLREFCLK_SEL  (3'b001),
            .SIM_VERSION         ("2.0"),


           //----------------COMMON BLOCK Attributes---------------
            .BIAS_CFG                               (64'h0000040000001050),
            .COMMON_CFG                             (32'h0000001C),
            .QPLL_CFG                               (27'h04801C7),
            .QPLL_CLKOUT_CFG                        (4'b1111),
            .QPLL_COARSE_FREQ_OVRD                  (6'b010000),
            .QPLL_COARSE_FREQ_OVRD_EN               (1'b0),
            .QPLL_CP                                (10'b0000011111),
            .QPLL_CP_MONITOR_EN                     (1'b0),
            .QPLL_DMONITOR_SEL                      (1'b0),
            .QPLL_FBDIV                             (QPLL_FBDIV_IN),
            .QPLL_FBDIV_MONITOR_EN                  (1'b0),
            .QPLL_FBDIV_RATIO                       (QPLL_FBDIV_RATIO),
            .QPLL_INIT_CFG                          (24'h000006),
            .QPLL_LOCK_CFG                          (16'h05E8),
            .QPLL_LPF                               (4'b1111),
            .QPLL_REFCLK_DIV                        (1),
            .RSVD_ATTR0                             (16'h0000),
            .RSVD_ATTR1                             (16'h0000),
            .QPLL_RP_COMP                           (1'b0),
            .QPLL_VTRL_RESET                        (2'b00),
            .RCAL_CFG                               (2'b00)

    )
    gthe2_common_0_i
    (
        //----------- Common Block  - Dynamic Reconfiguration Port (DRP) -----------
        .DRPADDR                        (tied_to_ground_vec_i[7:0]),
        .DRPCLK                         (tied_to_ground_i),
        .DRPDI                          (tied_to_ground_vec_i[15:0]),
        .DRPDO                          (),
        .DRPEN                          (tied_to_ground_i),
        .DRPRDY                         (),
        .DRPWE                          (tied_to_ground_i),
        //-------------------- Common Block  - Ref Clock Ports ---------------------
        .GTGREFCLK                      (GT0_GTGREFCLK_COMMON_IN),
        .GTNORTHREFCLK0                 (GT0_GTNORTHREFCLK0_COMMON_IN),
        .GTNORTHREFCLK1                 (GT0_GTNORTHREFCLK1_COMMON_IN),
        .GTREFCLK0                      (GT0_GTREFCLK0_COMMON_IN),
        .GTREFCLK1                      (GT0_GTREFCLK1_COMMON_IN),
        .GTSOUTHREFCLK0                 (GT0_GTSOUTHREFCLK0_COMMON_IN),
        .GTSOUTHREFCLK1                 (GT0_GTSOUTHREFCLK1_COMMON_IN),
        //----------------------- Common Block -  QPLL Ports -----------------------
        .QPLLDMONITOR                   (),
        //--------------------- Common Block - Clocking Ports ----------------------
        .QPLLOUTCLK                     (gt0_qplloutclk_i),
        .QPLLOUTREFCLK                  (gt0_qplloutrefclk_i),
        .REFCLKOUTMONITOR               (),
        //----------------------- Common Block - QPLL Ports ------------------------
        .BGRCALOVRDENB                  (tied_to_vcc_i),
        .PMARSVDOUT                     (),
        .QPLLFBCLKLOST                  (),
        .QPLLLOCK                       (GT0_QPLLLOCK_OUT),
        .QPLLLOCKDETCLK                 (GT0_QPLLLOCKDETCLK_IN),
        .QPLLLOCKEN                     (tied_to_vcc_i),
        .QPLLOUTRESET                   (tied_to_ground_i),
        .QPLLPD                         (tied_to_ground_i),
        .QPLLREFCLKLOST                 (GT0_QPLLREFCLKLOST_OUT),
        .QPLLREFCLKSEL                  (3'b001),
        .QPLLRESET                      (GT0_QPLLRESET_IN),
        .QPLLRSVD1                      (16'b0000000000000000),
        .QPLLRSVD2                      (5'b11111),
        //------------------------------- QPLL Ports -------------------------------
        .BGBYPASSB                      (tied_to_vcc_i),
        .BGMONITORENB                   (tied_to_vcc_i),
        .BGPDB                          (tied_to_vcc_i),
        .BGRCALOVRD                     (5'b00000),
        .PMARSVD                        (8'b00000000),
        .RCALENB                        (tied_to_vcc_i)

    );


endmodule

    
