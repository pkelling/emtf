//------------------------------------------------------------------------------
//   ____  ____
//  /   /\/   /
// /___/  \  /    Vendor: Xilinx
// \   \   \/     Version : 2.7
//  \   \         Application : 7 Series FPGAs Transceivers Wizard 
//  /   /         Filename : daq_link_tx_init.v
// /___/   /\      
// \   \  /  \ 
//  \___\/\___\
//
//  Description : This module instantiates the modules required for
//                reset and initialisation of the Transceiver
//
// Module daq_link_tx_init
// Generated by Xilinx 7 Series FPGAs Transceivers Wizard
// 
// 
// (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES. 


`timescale 1ns / 1ps
`define DLY #1

//***********************************Entity Declaration************************

module daq_link_tx_init #
(
    parameter EXAMPLE_SIM_GTRESET_SPEEDUP            = "TRUE",                  // Simulation setting for GT SecureIP model
    parameter EXAMPLE_SIMULATION                     =  0,                      // Set to 1 for simulation
    parameter STABLE_CLOCK_PERIOD                    =  16, // Period of the stable clock driving this 
                                                                                // state-machine, unit is [ns]

    parameter EXAMPLE_USE_CHIPSCOPE                  =  0                       // Set to 1 to use Chipscope to drive resets

)
(
    input           SYSCLK_IN,
    input           SOFT_RESET_IN,
    input           DONT_RESET_ON_DATA_ERROR_IN,
    output          GT0_TX_FSM_RESET_DONE_OUT,
    output          GT0_RX_FSM_RESET_DONE_OUT,
    input           GT0_DATA_VALID_IN,

    //_________________________________________________________________________
    //GT0  (X0Y0)
    //____________________________CHANNEL PORTS________________________________
    //------------------------------- CPLL Ports -------------------------------
    output          GT0_CPLLFBCLKLOST_OUT,
    output          GT0_CPLLLOCK_OUT,
    input           GT0_CPLLLOCKDETCLK_IN,
    input           GT0_CPLLRESET_IN,
    //------------------------ Channel - Clocking Ports ------------------------
    input           GT0_GTREFCLK0_IN,
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   GT0_DRPADDR_IN,
    input           GT0_DRPCLK_IN,
    input   [15:0]  GT0_DRPDI_IN,
    output  [15:0]  GT0_DRPDO_OUT,
    input           GT0_DRPEN_IN,
    output          GT0_DRPRDY_OUT,
    input           GT0_DRPWE_IN,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          GT0_EYESCANDATAERROR_OUT,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           GT0_GTRXRESET_IN,
    //------------------- TX Initialization and Reset Ports --------------------
    input           GT0_GTTXRESET_IN,
    input           GT0_TXUSERRDY_IN,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           GT0_TXUSRCLK_IN,
    input           GT0_TXUSRCLK2_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [15:0]  GT0_TXDATA_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GT0_GTHTXN_OUT,
    output          GT0_GTHTXP_OUT,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          GT0_TXOUTCLK_OUT,
    output          GT0_TXOUTCLKFABRIC_OUT,
    output          GT0_TXOUTCLKPCS_OUT,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          GT0_TXRESETDONE_OUT,
    //--------------- Transmit Ports - TX Polarity Control Ports ---------------
    input           GT0_TXPOLARITY_IN,
    //---------------- Transmit Ports - pattern Generator Ports ----------------
    input   [2:0]   GT0_TXPRBSSEL_IN,
    //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    input   [1:0]   GT0_TXCHARISK_IN,


    //____________________________COMMON PORTS________________________________
    //-------------------- Common Block  - Ref Clock Ports ---------------------
    input           GT0_GTREFCLK0_COMMON_IN,
    //----------------------- Common Block - QPLL Ports ------------------------
    output          GT0_QPLLLOCK_OUT,
    input           GT0_QPLLLOCKDETCLK_IN,
    input           GT0_QPLLRESET_IN


);



//***********************************Parameter Declarations********************

    //Typical CDRLOCK Time is 50,000UI, as per DS183
    localparam RX_CDRLOCK_TIME      = (EXAMPLE_SIMULATION == 1) ? 1000 : 50000/5;

       
    integer   WAIT_TIME_CDRLOCK    = RX_CDRLOCK_TIME / STABLE_CLOCK_PERIOD;      

//-------------------------- GT Wrapper Wires ------------------------------
    wire           gt0_cpllreset_i;
    wire           gt0_cpllreset_t;
    wire           gt0_cpllrefclklost_i;
    wire           gt0_cplllock_i;
    wire           gt0_txresetdone_i;
    wire           gt0_rxresetdone_i;
    wire           gt0_gttxreset_i;
    wire           gt0_gttxreset_t;
    wire           gt0_gtrxreset_i;
    wire           gt0_gtrxreset_t;
    wire           gt0_txuserrdy_i;
    wire           gt0_txuserrdy_t;
    wire           gt0_rxuserrdy_i;
    wire           gt0_rxuserrdy_t;

    wire           gt0_rxdfeagchold_i;
    wire           gt0_rxdfelfhold_i;
    wire           gt0_rxlpmlfhold_i;
    wire           gt0_rxlpmhfhold_i;



    wire           gt0_qpllreset_i;
    wire           gt0_qpllreset_t;
    wire           gt0_qpllrefclklost_i;
    wire           gt0_qplllock_i;


//------------------------------- Global Signals -----------------------------
    wire           tied_to_ground_i;
    wire           tied_to_vcc_i;










 


//**************************** Main Body of Code *******************************
    //  Static signal Assigments
    assign  tied_to_ground_i                     =  1'b0;
    assign  tied_to_vcc_i                        =  1'b1;

//    ----------------------------- The GT Wrapper -----------------------------
    
    // Use the instantiation template in the example directory to add the GT wrapper to your design.
    // In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    // checker. The GTs will reset, then attempt to align and transmit data. If channel bonding is 
    // enabled, bonding should occur after alignment.


    daq_link_tx #
    (
        .EXAMPLE_SIMULATION             (EXAMPLE_SIMULATION),
        .WRAPPER_SIM_GTRESET_SPEEDUP    (EXAMPLE_SIM_GTRESET_SPEEDUP)
    )
    daq_link_tx_i
    (
  
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT0  (X0Y0)

        //------------------------------- CPLL Ports -------------------------------
        .GT0_CPLLFBCLKLOST_OUT          (GT0_CPLLFBCLKLOST_OUT),
        .GT0_CPLLLOCK_OUT               (gt0_cplllock_i),
        .GT0_CPLLLOCKDETCLK_IN          (GT0_CPLLLOCKDETCLK_IN),
        .GT0_CPLLREFCLKLOST_OUT         (gt0_cpllrefclklost_i),
        .GT0_CPLLRESET_IN               (gt0_cpllreset_i),
        //------------------------ Channel - Clocking Ports ------------------------
        .GT0_GTREFCLK0_IN               (GT0_GTREFCLK0_IN),
        //-------------------------- Channel - DRP Ports  --------------------------
        .GT0_DRPADDR_IN                 (GT0_DRPADDR_IN),
        .GT0_DRPCLK_IN                  (GT0_DRPCLK_IN),
        .GT0_DRPDI_IN                   (GT0_DRPDI_IN),
        .GT0_DRPDO_OUT                  (GT0_DRPDO_OUT),
        .GT0_DRPEN_IN                   (GT0_DRPEN_IN),
        .GT0_DRPRDY_OUT                 (GT0_DRPRDY_OUT),
        .GT0_DRPWE_IN                   (GT0_DRPWE_IN),
        //------------------------ RX Margin Analysis Ports ------------------------
        .GT0_EYESCANDATAERROR_OUT       (GT0_EYESCANDATAERROR_OUT),
        //------------------- Receive Ports - RX Equalizer Ports -------------------
        .GT0_RXDFEAGCHOLD_IN            (gt0_rxdfeagchold_i),
        .GT0_RXDFELFHOLD_IN             (gt0_rxdfelfhold_i),
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .GT0_GTRXRESET_IN               (gt0_gtrxreset_i),
        //------------------- TX Initialization and Reset Ports --------------------
        .GT0_GTTXRESET_IN               (gt0_gttxreset_i),
        .GT0_TXUSERRDY_IN               (gt0_txuserrdy_i),
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .GT0_TXUSRCLK_IN                (GT0_TXUSRCLK_IN),
        .GT0_TXUSRCLK2_IN               (GT0_TXUSRCLK2_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GT0_TXDATA_IN                  (GT0_TXDATA_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GT0_GTHTXN_OUT                 (GT0_GTHTXN_OUT),
        .GT0_GTHTXP_OUT                 (GT0_GTHTXP_OUT),
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .GT0_TXOUTCLK_OUT               (GT0_TXOUTCLK_OUT),
        .GT0_TXOUTCLKFABRIC_OUT         (GT0_TXOUTCLKFABRIC_OUT),
        .GT0_TXOUTCLKPCS_OUT            (GT0_TXOUTCLKPCS_OUT),
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .GT0_TXRESETDONE_OUT            (gt0_txresetdone_i),
        //--------------- Transmit Ports - TX Polarity Control Ports ---------------
        .GT0_TXPOLARITY_IN              (GT0_TXPOLARITY_IN),
        //---------------- Transmit Ports - pattern Generator Ports ----------------
        .GT0_TXPRBSSEL_IN               (GT0_TXPRBSSEL_IN),
        //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        .GT0_TXCHARISK_IN               (GT0_TXCHARISK_IN),




    //____________________________COMMON PORTS________________________________
        //-------------------- Common Block  - Ref Clock Ports ---------------------
        .GT0_GTREFCLK0_COMMON_IN        (GT0_GTREFCLK0_COMMON_IN),
        //----------------------- Common Block - QPLL Ports ------------------------
        .GT0_QPLLLOCK_OUT               (gt0_qplllock_i),
        .GT0_QPLLLOCKDETCLK_IN          (GT0_QPLLLOCKDETCLK_IN),
        .GT0_QPLLREFCLKLOST_OUT         (gt0_qpllrefclklost_i),
        .GT0_QPLLRESET_IN               (gt0_qpllreset_i)

    );




    assign  GT0_CPLLLOCK_OUT                     =  gt0_cplllock_i;
    assign  GT0_TXRESETDONE_OUT                  =  gt0_txresetdone_i;
    assign  GT0_QPLLLOCK_OUT                     =  gt0_qplllock_i;

generate
if (EXAMPLE_USE_CHIPSCOPE == 1) 
begin : chipscope
    assign  gt0_cpllreset_i                      =  GT0_CPLLRESET_IN || gt0_cpllreset_t;
    assign  gt0_gttxreset_i                      =  GT0_GTTXRESET_IN || gt0_gttxreset_t;
    assign  gt0_gtrxreset_i                      =  GT0_GTRXRESET_IN || gt0_gtrxreset_t;
    assign  gt0_txuserrdy_i                      =  GT0_TXUSERRDY_IN || gt0_txuserrdy_t;
    assign  gt0_qpllreset_i                      =  GT0_QPLLRESET_IN || gt0_qpllreset_t;
end
endgenerate 

generate
if (EXAMPLE_USE_CHIPSCOPE == 0) 
begin : no_chipscope
    assign  gt0_cpllreset_i                      =  gt0_cpllreset_t;
    assign  gt0_gttxreset_i                      =  gt0_gttxreset_t;
    assign  gt0_gtrxreset_i                      =  gt0_gtrxreset_t;
    assign  gt0_txuserrdy_i                      =  gt0_txuserrdy_t;
    assign  gt0_rxuserrdy_i                      =  gt0_rxuserrdy_t;
    assign  gt0_qpllreset_i                      =  gt0_qpllreset_t;
end
endgenerate 


daq_link_tx_TX_STARTUP_FSM #
          (
           .GT_TYPE                  ("GTH"), //GTX or GTH or GTP
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("FALSE"),                       // the TX and RX Reset FSMs must
           .RX_QPLL_USED             ("FALSE"),                       // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt0_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (SYSCLK_IN),
        .TXUSERCLK                      (GT0_TXUSRCLK_IN),
        .SOFT_RESET                     (SOFT_RESET_IN),
        .QPLLREFCLKLOST                 (tied_to_ground_i),
        .CPLLREFCLKLOST                 (gt0_cpllrefclklost_i),
        .QPLLLOCK                       (tied_to_vcc_i),
        .CPLLLOCK                       (gt0_cplllock_i),
        .TXRESETDONE                    (gt0_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt0_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (gt0_cpllreset_t),
        .TX_FSM_RESET_DONE              (GT0_TX_FSM_RESET_DONE_OUT),
        .TXUSERRDY                      (gt0_txuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RETRY_COUNTER                  ()
           );











endmodule


